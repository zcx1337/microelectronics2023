library verilog;
use verilog.vl_types.all;
entity TIMER_tb is
end TIMER_tb;
